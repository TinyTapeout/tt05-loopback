/*
 * tt_um_loopback.v
 *
 * Loopback test user module
 *
 * Author: Sylvain Munaut <tnt@246tNt.com>
 */

`default_nettype none

module tt_um_loopback (
	input  wire [7:0] ui_in,	// Dedicated inputs
	output wire [7:0] uo_out,	// Dedicated outputs
	input  wire [7:0] uio_in,	// IOs: Input path
	output wire [7:0] uio_out,	// IOs: Output path
	output wire [7:0] uio_oe,	// IOs: Enable path (active high: 0=input, 1=output)
	input  wire       ena,
	input  wire       clk,
	input  wire       rst_n
);

	assign uo_out[6:0] = {7{ui_in[0]}};
	assign uo_out[7] = &ui_in[7:4];

	assign uio_out = 0;
	assign uio_oe = 0;

endmodule // tt_um_loopback
